module toUpper (in,out);
    input [7:0] in; 
    output [7:0] out;
    wire a0, a1, a2, a3, a4, a5, a6, a7;

    
  
    
endmodule